
module arb # (
) (

);

// fairly choose 1 or 2 (depending on output buses) cmds
// mark taken from queue
// obey restrictions from smp, etc.
// detect addr collisions - not needed if no caching?


endmodule